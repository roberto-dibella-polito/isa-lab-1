-- Project 1: IIR filter
-- Constants

package constants is

	constant numBit : integer := 8;
	
end constants;